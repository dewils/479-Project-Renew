magic
tech scmos
timestamp 1428875432
<< pwell >>
rect 2 18 14 35
<< nwell >>
rect 2 35 14 48
<< polysilicon >>
rect 7 48 9 50
rect 7 30 9 40
rect 7 24 9 26
<< ndiffusion >>
rect 6 26 7 30
rect 9 26 10 30
<< pdiffusion >>
rect 6 40 7 48
rect 9 40 10 48
<< metal1 >>
rect 2 56 6 65
rect 2 52 10 56
rect 2 48 6 52
rect 11 37 14 40
rect 2 33 3 37
rect 11 30 14 33
rect 2 22 6 26
rect 2 18 10 22
rect 2 9 6 18
<< metal2 >>
rect -6 65 2 69
rect 6 65 19 69
rect -6 34 -2 37
rect 15 33 19 36
rect -6 5 2 9
rect 6 5 19 9
<< ntransistor >>
rect 7 26 9 30
<< ptransistor >>
rect 7 40 9 48
<< polycontact >>
rect 3 33 7 37
<< ndcontact >>
rect 2 26 6 30
rect 10 26 14 30
<< pdcontact >>
rect 2 40 6 48
rect 10 40 14 48
<< m2contact >>
rect 2 65 6 69
rect -2 33 2 37
rect 11 33 15 37
rect 2 5 6 9
<< psubstratepcontact >>
rect 10 18 14 22
<< nsubstratencontact >>
rect 10 52 14 56
<< labels >>
rlabel metal2 15 33 19 36 3 Y
rlabel metal2 6 65 19 69 3 Vdd
rlabel metal2 6 5 19 9 3 GND
rlabel metal2 -6 65 2 69 7 Vdd
rlabel metal2 -6 5 2 9 7 GND
rlabel metal2 -6 34 -2 37 7 A
<< end >>
