magic
tech scmos
timestamp 1428895890
<< metal1 >>
rect -12 922 -8 986
rect -12 822 -8 918
rect -12 709 -8 818
rect -12 596 -8 705
rect -12 483 -8 592
rect -12 370 -8 479
rect -12 257 -8 366
rect -12 144 -8 253
rect -12 31 -8 140
rect -12 -8 -8 27
rect -12 -16 -8 -12
rect -4 982 0 986
rect -4 882 0 978
rect 15 950 18 986
rect 127 950 130 986
rect 178 950 181 986
rect 15 904 18 946
rect 43 908 46 945
rect 127 908 130 946
rect 155 904 158 946
rect 178 904 181 946
rect 192 904 195 986
rect 288 951 291 986
rect 220 908 223 946
rect 288 904 291 947
rect 316 908 319 946
rect 471 904 474 986
rect 486 922 490 986
rect -4 769 0 878
rect -4 656 0 765
rect -4 543 0 652
rect -4 430 0 539
rect -4 317 0 426
rect -4 204 0 313
rect -4 91 0 200
rect -4 0 0 87
rect 486 822 490 918
rect 486 709 490 818
rect 486 596 490 705
rect 486 483 490 592
rect 486 370 490 479
rect 486 257 490 366
rect 486 144 490 253
rect 486 31 490 140
rect -4 -16 0 -4
rect 192 -16 195 0
rect 486 -8 490 27
rect 486 -16 490 -12
rect 494 982 498 986
rect 494 882 498 978
rect 494 769 498 878
rect 494 656 498 765
rect 494 543 498 652
rect 494 430 498 539
rect 494 317 498 426
rect 494 204 498 313
rect 494 91 498 200
rect 494 0 498 87
rect 494 -16 498 -4
<< metal2 >>
rect 0 978 18 982
rect 43 978 130 982
rect 146 978 195 982
rect 199 978 291 982
rect 316 978 494 982
rect 182 947 195 950
rect -8 918 18 922
rect 43 918 130 922
rect 146 918 195 922
rect 199 918 291 922
rect 316 918 486 922
rect 26 904 42 907
rect 131 904 147 907
rect 189 904 219 907
rect 285 904 315 907
rect 486 878 494 882
rect -16 856 0 859
rect 486 845 502 848
rect -8 818 0 822
rect 486 765 494 769
rect -16 743 0 746
rect 486 732 502 735
rect -8 705 0 709
rect 486 652 494 656
rect -16 630 0 633
rect 486 619 502 622
rect -8 592 0 596
rect 486 539 494 543
rect -16 517 0 520
rect 486 506 502 509
rect -8 479 0 483
rect 486 426 494 430
rect -16 404 0 407
rect 486 393 502 396
rect -8 366 0 370
rect 486 313 494 317
rect -16 291 0 294
rect 486 280 502 283
rect -8 253 0 257
rect 486 200 494 204
rect -16 178 0 181
rect 486 167 502 170
rect -8 140 0 144
rect 486 87 494 91
rect -16 65 0 68
rect 486 54 502 57
rect -8 27 0 31
rect -16 -4 -4 0
rect 0 -4 494 0
rect 498 -4 502 0
rect -16 -12 -12 -8
rect -8 -12 486 -8
rect 490 -12 502 -8
<< m2contact >>
rect -12 918 -8 922
rect -12 818 -8 822
rect -12 705 -8 709
rect -12 592 -8 596
rect -12 479 -8 483
rect -12 366 -8 370
rect -12 253 -8 257
rect -12 140 -8 144
rect -12 27 -8 31
rect -12 -12 -8 -8
rect -4 978 0 982
rect 14 946 18 950
rect 42 945 46 949
rect 126 946 130 950
rect 22 904 26 908
rect 42 904 46 908
rect 155 946 159 950
rect 178 946 182 950
rect 127 904 131 908
rect 147 904 151 908
rect 185 904 189 908
rect 220 946 224 950
rect 287 947 291 951
rect 219 904 223 908
rect 281 904 285 908
rect 316 946 320 950
rect 315 904 319 908
rect 486 918 490 922
rect -4 878 0 882
rect -4 765 0 769
rect -4 652 0 656
rect -4 539 0 543
rect -4 426 0 430
rect -4 313 0 317
rect -4 200 0 204
rect -4 87 0 91
rect 486 818 490 822
rect 486 705 490 709
rect 486 592 490 596
rect 486 479 490 483
rect 486 366 490 370
rect 486 253 490 257
rect 486 140 490 144
rect 486 27 490 31
rect -4 -4 0 0
rect 486 -12 490 -8
rect 494 978 498 982
rect 494 878 498 882
rect 494 765 498 769
rect 494 652 498 656
rect 494 539 498 543
rect 494 426 498 430
rect 494 313 498 317
rect 494 200 498 204
rect 494 87 498 91
rect 494 -4 498 0
use ../cells/inverter1  inverter1_0
timestamp 1428875432
transform 1 0 24 0 1 913
box -6 5 19 69
use ../cells/inverter1  inverter1_1
timestamp 1428875432
transform 1 0 136 0 1 913
box -6 5 19 69
use ../cells/inverter1  inverter1_2
timestamp 1428875432
transform 1 0 201 0 1 913
box -6 5 19 69
use ../cells/inverter1  inverter1_3
timestamp 1428875432
transform 1 0 297 0 1 913
box -6 5 19 69
use dbitlow  dbitlow_0
array 0 0 486 0 7 113
timestamp 1428883144
transform 1 0 19 0 1 36
box -19 -36 467 77
<< labels >>
rlabel metal1 -12 922 -8 986 1 GND
rlabel metal1 -4 982 0 986 1 Vdd
rlabel metal1 494 982 498 986 1 Vdd
rlabel metal1 486 922 490 986 1 GND
rlabel metal1 15 950 18 986 1 S0
rlabel metal1 127 950 130 986 1 S1
rlabel metal1 178 950 181 986 1 shift
rlabel metal1 192 904 195 986 1 inbit
rlabel metal1 288 951 291 986 1 clk
rlabel metal1 471 904 474 986 1 reset_n
rlabel metal2 486 845 502 848 3 quotient_0
rlabel metal2 486 732 502 735 3 quotient_1
rlabel metal2 486 619 502 622 3 quotient_2
rlabel metal2 486 506 502 509 3 quotient_3
rlabel metal2 486 393 502 396 3 quotient_4
rlabel metal2 486 280 502 283 3 quotient_5
rlabel metal2 486 167 502 170 3 quotient_6
rlabel metal2 486 54 502 57 3 quotient_7
rlabel metal1 192 -16 195 0 5 outbit
rlabel metal1 -4 -16 0 -4 5 Vdd
rlabel metal1 -12 -16 -8 -12 5 GND
rlabel metal2 -16 65 0 68 7 dividendin_7
rlabel metal2 -16 178 0 181 7 dividendin_6
rlabel metal2 -16 291 0 294 7 dividendin_5
rlabel metal2 -16 404 0 407 7 dividendin_4
rlabel metal2 -16 517 0 520 7 dividendin_3
rlabel metal2 -16 630 0 633 7 dividendin_2
rlabel metal2 -16 743 0 746 7 dividendin_1
rlabel metal2 -16 856 0 859 7 dividendin_0
rlabel metal1 494 -16 498 -4 5 Vdd
rlabel metal1 486 -16 490 -12 5 GND
<< end >>
