magic
tech scmos
timestamp 1428902219
<< pwell >>
rect -1 3 61 24
<< nwell >>
rect -1 24 61 49
<< polysilicon >>
rect 4 15 6 56
rect 20 15 22 56
rect 38 41 40 43
rect 54 41 56 43
rect 38 15 40 33
rect 54 15 56 33
rect 4 9 6 11
rect 20 9 22 11
rect 38 9 40 11
rect 54 9 56 11
<< ndiffusion >>
rect 3 11 4 15
rect 6 11 7 15
rect 19 11 20 15
rect 22 11 23 15
rect 37 11 38 15
rect 40 11 41 15
rect 53 11 54 15
rect 56 11 57 15
<< pdiffusion >>
rect 37 33 38 41
rect 40 33 41 41
rect 53 33 54 41
rect 56 33 57 41
<< metal1 >>
rect -22 74 -19 77
rect -22 -23 -19 70
rect -15 67 -12 77
rect -15 -23 -12 63
rect -8 28 -5 77
rect 7 56 10 63
rect 23 56 26 70
rect -1 49 3 55
rect 57 49 61 55
rect -1 45 33 49
rect 37 45 49 49
rect 53 45 61 49
rect 33 41 37 45
rect 49 41 53 45
rect -8 -23 -5 16
rect -1 15 2 16
rect 8 15 11 16
rect 15 15 18 24
rect 42 25 45 33
rect 58 25 61 33
rect 34 21 37 25
rect 28 18 37 21
rect 42 21 50 25
rect 24 15 27 17
rect 42 15 45 21
rect 58 15 61 21
rect 33 7 37 11
rect 49 7 53 11
rect -1 3 11 7
rect 15 3 33 7
rect 37 3 49 7
rect 53 3 61 7
rect -1 -1 3 3
rect 57 -1 61 3
<< metal2 >>
rect -19 71 22 74
rect -11 63 7 66
rect -26 55 -1 59
rect 61 55 73 59
rect -5 24 14 27
rect 62 22 73 25
rect -26 16 -9 19
rect -5 16 -2 20
rect 12 17 24 20
rect -26 -5 -1 -1
rect 61 -5 73 -1
<< ntransistor >>
rect 4 11 6 15
rect 20 11 22 15
rect 38 11 40 15
rect 54 11 56 15
<< ptransistor >>
rect 38 33 40 41
rect 54 33 56 41
<< polycontact >>
rect 6 52 10 56
rect 22 52 26 56
rect 34 25 38 29
rect 50 21 54 25
<< ndcontact >>
rect -1 11 3 15
rect 7 11 11 15
rect 15 11 19 15
rect 23 11 27 15
rect 33 11 37 15
rect 41 11 45 15
rect 49 11 53 15
rect 57 11 61 15
<< pdcontact >>
rect 33 33 37 41
rect 41 33 45 41
rect 49 33 53 41
rect 57 33 61 41
<< m2contact >>
rect -23 70 -19 74
rect -15 63 -11 67
rect 22 70 26 74
rect 7 63 11 67
rect -1 55 3 59
rect 57 55 61 59
rect -9 24 -5 28
rect 14 24 18 28
rect -9 16 -5 20
rect -2 16 2 20
rect 8 16 12 20
rect 24 17 28 21
rect 58 21 62 25
rect -1 -5 3 -1
rect 57 -5 61 -1
<< psubstratepcontact >>
rect 11 3 15 7
rect 33 3 37 7
rect 49 3 53 7
<< nsubstratencontact >>
rect 33 45 37 49
rect 49 45 53 49
<< labels >>
rlabel metal1 -22 74 -19 77 1 shift
rlabel metal1 -15 67 -12 77 1 shift_n
rlabel metal1 -8 28 -5 77 1 inbit
rlabel metal2 -26 55 -1 59 7 Vdd
rlabel metal2 -26 16 -9 19 7 A
rlabel metal2 -26 -5 -1 -1 7 GND
rlabel metal1 -22 -23 -19 70 5 shift
rlabel metal1 -15 -23 -12 63 5 shift_n
rlabel metal1 -8 -23 -5 16 5 A
rlabel metal2 61 55 73 59 3 Vdd
rlabel metal2 62 22 73 25 3 B
rlabel metal2 61 -5 73 -1 3 GND
<< end >>
