magic
tech scmos
timestamp 1428878105
<< pwell >>
rect -55 28 12 50
<< nwell >>
rect -55 50 12 79
<< polysilicon >>
rect -50 71 -48 87
rect -34 71 -32 82
rect -16 71 -14 87
rect 1 71 3 82
rect -50 52 -48 63
rect -34 59 -32 63
rect -34 57 -23 59
rect -50 50 -32 52
rect -50 40 -48 42
rect -34 40 -32 50
rect -50 27 -48 36
rect -34 34 -32 36
rect -25 27 -23 57
rect -16 48 -14 63
rect 1 56 3 63
rect 1 54 12 56
rect -16 46 3 48
rect -16 40 -14 42
rect 1 40 3 46
rect -50 25 -23 27
rect -16 27 -14 36
rect 1 34 3 36
rect 10 27 12 54
rect -16 25 12 27
<< ndiffusion >>
rect -51 36 -50 40
rect -48 36 -47 40
rect -35 36 -34 40
rect -32 36 -31 40
rect -17 36 -16 40
rect -14 36 -13 40
rect 0 36 1 40
rect 3 36 4 40
<< pdiffusion >>
rect -51 63 -50 71
rect -48 63 -47 71
rect -35 63 -34 71
rect -32 63 -31 71
rect -17 63 -16 71
rect -14 63 -13 71
rect 0 63 1 71
rect 3 63 4 71
<< metal1 >>
rect -83 92 -80 102
rect -83 3 -80 88
rect -76 99 -73 102
rect -76 3 -73 95
rect -47 87 -46 91
rect -34 86 -31 94
rect -18 87 -17 91
rect 0 86 3 95
rect 16 92 19 102
rect 23 100 26 102
rect -55 79 -51 80
rect 8 79 12 80
rect -55 75 -43 79
rect -39 75 -26 79
rect -22 75 -9 79
rect -5 75 12 79
rect -55 61 -52 63
rect -69 16 -66 49
rect -62 8 -59 41
rect -55 40 -52 57
rect -46 61 -43 63
rect -46 40 -43 57
rect -39 46 -36 63
rect -39 40 -36 42
rect -30 46 -27 63
rect -21 61 -18 63
rect -21 45 -18 57
rect -30 40 -27 42
rect -21 40 -18 41
rect -12 61 -9 63
rect -12 40 -9 57
rect -4 53 -1 63
rect 5 62 8 63
rect 5 53 8 58
rect -4 40 -1 49
rect 5 40 8 49
rect -55 28 -43 32
rect -39 28 -22 32
rect -18 28 -9 32
rect -5 28 12 32
rect -55 24 -51 28
rect 8 24 12 28
rect 16 2 19 88
rect 23 2 26 96
<< metal2 >>
rect -72 95 -35 98
rect 4 96 23 99
rect -80 88 -46 91
rect -18 88 16 91
rect -87 80 -55 84
rect 12 80 30 84
rect -87 57 -56 60
rect -42 57 -22 60
rect -8 58 5 61
rect -87 50 -70 53
rect -66 50 -4 53
rect 9 50 30 53
rect -87 42 -63 45
rect -59 42 -40 45
rect -26 42 -22 45
rect -87 20 -55 24
rect 12 20 30 24
rect -66 13 30 16
rect -59 5 30 8
<< ntransistor >>
rect -50 36 -48 40
rect -34 36 -32 40
rect -16 36 -14 40
rect 1 36 3 40
<< ptransistor >>
rect -50 63 -48 71
rect -34 63 -32 71
rect -16 63 -14 71
rect 1 63 3 71
<< polycontact >>
rect -51 87 -47 91
rect -17 87 -13 91
rect -35 82 -31 86
rect 0 82 4 86
<< ndcontact >>
rect -55 36 -51 40
rect -47 36 -43 40
rect -39 36 -35 40
rect -31 36 -27 40
rect -43 28 -39 32
rect -21 36 -17 40
rect -13 36 -9 40
rect -4 36 0 40
rect 4 36 8 40
rect -22 28 -18 32
rect -9 28 -5 32
<< pdcontact >>
rect -43 75 -39 79
rect -26 75 -22 79
rect -9 75 -5 79
rect -55 63 -51 71
rect -47 63 -43 71
rect -39 63 -35 71
rect -31 63 -27 71
rect -21 63 -17 71
rect -13 63 -9 71
rect -4 63 0 71
rect 4 63 8 71
<< m2contact >>
rect -84 88 -80 92
rect -76 95 -72 99
rect -35 94 -31 98
rect -46 87 -42 91
rect 0 95 4 99
rect -22 87 -18 91
rect -55 80 -51 84
rect 23 96 27 100
rect 16 88 20 92
rect 8 80 12 84
rect -56 57 -52 61
rect -70 49 -66 53
rect -63 41 -59 45
rect -70 12 -66 16
rect -46 57 -42 61
rect -40 42 -36 46
rect -22 57 -18 61
rect -30 42 -26 46
rect -22 41 -18 45
rect -12 57 -8 61
rect 5 58 9 62
rect -4 49 0 53
rect 5 49 9 53
rect -55 20 -51 24
rect 8 20 12 24
rect -63 4 -59 8
<< labels >>
rlabel metal1 -83 3 -80 88 5 S0
rlabel metal1 -76 3 -73 95 5 S0_n
rlabel metal1 16 92 19 102 1 S1
rlabel metal1 23 100 26 102 1 S1_n
rlabel metal1 16 2 19 88 5 S1
rlabel metal1 23 2 26 96 5 S1_n
rlabel metal2 -87 80 -55 84 7 Vdd
rlabel metal2 -87 20 -55 24 7 GND
rlabel metal2 12 80 30 84 3 Vdd
rlabel metal2 12 20 30 24 3 GND
rlabel metal2 -87 57 -56 60 7 D0
rlabel metal2 -87 50 -70 53 7 D1
rlabel metal2 -87 42 -63 45 7 D2
rlabel metal2 -66 13 30 16 3 D1
rlabel metal2 -59 5 30 8 3 D2
rlabel metal1 -83 92 -80 102 1 S0
rlabel metal1 -76 99 -73 102 1 S0_n
rlabel metal2 9 50 30 53 3 Y
<< end >>
