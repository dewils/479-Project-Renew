magic
tech scmos
timestamp 1428289220
<< pwell >>
rect -58 28 61 50
<< nwell >>
rect -58 50 61 77
<< polysilicon >>
rect -49 69 -47 100
rect -33 69 -31 100
rect -17 69 -15 71
rect 0 69 2 71
rect 17 69 19 100
rect 33 69 35 100
rect 49 69 51 71
rect -49 59 -47 61
rect -33 59 -31 61
rect -17 46 -15 61
rect 0 58 2 61
rect 17 59 19 61
rect 33 59 35 61
rect 49 57 51 61
rect 44 55 51 57
rect -22 44 -15 46
rect -49 40 -47 42
rect -33 40 -31 42
rect -17 40 -15 44
rect 0 40 2 44
rect 17 40 19 42
rect 33 40 35 42
rect 49 40 51 55
rect -49 0 -47 36
rect -33 0 -31 36
rect -17 34 -15 36
rect 0 34 2 36
rect 17 0 19 36
rect 33 0 35 36
rect 49 34 51 36
<< ndiffusion >>
rect -50 36 -49 40
rect -47 36 -46 40
rect -34 36 -33 40
rect -31 36 -30 40
rect -18 36 -17 40
rect -15 36 -13 40
rect -1 36 0 40
rect 2 36 4 40
rect 16 36 17 40
rect 19 36 20 40
rect 32 36 33 40
rect 35 36 36 40
rect 48 36 49 40
rect 51 36 53 40
<< pdiffusion >>
rect -50 61 -49 69
rect -47 61 -46 69
rect -34 61 -33 69
rect -31 61 -30 69
rect -18 61 -17 69
rect -15 61 -13 69
rect -1 61 0 69
rect 2 61 4 69
rect 16 61 17 69
rect 19 61 20 69
rect 32 61 33 69
rect 35 61 36 69
rect 48 61 49 69
rect 51 61 53 69
<< metal1 >>
rect -58 73 -42 77
rect -38 73 -18 77
rect -14 73 -1 77
rect 3 73 24 77
rect 28 73 44 77
rect 48 73 61 77
rect -22 69 -18 73
rect -5 69 -1 73
rect 44 69 48 73
rect -54 60 -51 61
rect -54 40 -51 56
rect -45 60 -42 61
rect -45 40 -42 56
rect -38 45 -35 61
rect -38 40 -35 41
rect -29 60 -26 61
rect -29 40 -26 56
rect -12 45 -9 61
rect 5 60 8 61
rect -2 53 1 54
rect -2 48 1 49
rect -12 40 -9 41
rect 5 40 8 56
rect 12 45 15 61
rect 12 40 15 41
rect 21 45 24 61
rect 28 60 31 61
rect 21 40 24 41
rect 28 40 31 56
rect 37 45 40 61
rect 54 52 57 61
rect 37 40 40 41
rect 54 40 57 48
rect -22 32 -18 36
rect -5 32 -1 36
rect 44 32 48 36
rect -58 28 -42 32
rect -38 28 -19 32
rect -15 28 -1 32
rect 3 28 24 32
rect 28 28 44 32
rect 48 28 61 32
<< metal2 >>
rect -58 56 -55 59
rect -41 56 -29 59
rect 9 56 27 59
rect -58 49 -3 52
rect 58 49 61 52
rect -58 42 -39 45
rect -8 41 11 44
rect 25 41 37 44
<< ntransistor >>
rect -49 36 -47 40
rect -33 36 -31 40
rect -17 36 -15 40
rect 0 36 2 40
rect 17 36 19 40
rect 33 36 35 40
rect 49 36 51 40
<< ptransistor >>
rect -49 61 -47 69
rect -33 61 -31 69
rect -17 61 -15 69
rect 0 61 2 69
rect 17 61 19 69
rect 33 61 35 69
rect 49 61 51 69
<< polycontact >>
rect -26 43 -22 47
rect -2 54 2 58
rect 40 54 44 58
rect -2 44 2 48
<< ndcontact >>
rect -54 36 -50 40
rect -46 36 -42 40
rect -38 36 -34 40
rect -30 36 -26 40
rect -22 36 -18 40
rect -13 36 -9 40
rect -5 36 -1 40
rect 4 36 8 40
rect 12 36 16 40
rect 20 36 24 40
rect 28 36 32 40
rect 36 36 40 40
rect 44 36 48 40
rect 53 36 57 40
rect -42 28 -38 32
rect -19 28 -15 32
rect -1 28 3 32
rect 24 28 28 32
rect 44 28 48 32
<< pdcontact >>
rect -42 73 -38 77
rect -18 73 -14 77
rect -1 73 3 77
rect 24 73 28 77
rect 44 73 48 77
rect -54 61 -50 69
rect -46 61 -42 69
rect -38 61 -34 69
rect -30 61 -26 69
rect -22 61 -18 69
rect -13 61 -9 69
rect -5 61 -1 69
rect 4 61 8 69
rect 12 61 16 69
rect 20 61 24 69
rect 28 61 32 69
rect 36 61 40 69
rect 44 61 48 69
rect 53 61 57 69
<< m2contact >>
rect -55 56 -51 60
rect -45 56 -41 60
rect -39 41 -35 45
rect -29 56 -25 60
rect 5 56 9 60
rect -3 49 1 53
rect -12 41 -8 45
rect 11 41 15 45
rect 27 56 31 60
rect 21 41 25 45
rect 54 48 58 52
rect 37 41 41 45
<< labels >>
rlabel metal2 -58 56 -55 59 7 D0
rlabel metal2 -58 49 -3 52 7 D1
rlabel metal2 -58 42 -39 45 7 D2
rlabel metal2 58 49 61 52 3 Y
rlabel polysilicon -49 69 -47 100 1 S0
rlabel polysilicon -33 69 -31 100 1 S0_n
rlabel polysilicon 17 69 19 100 1 S1
rlabel polysilicon 33 69 35 100 1 S1_n
rlabel polysilicon -49 0 -47 36 5 S0_n
rlabel polysilicon -33 0 -31 36 5 S0
rlabel polysilicon 17 0 19 36 5 S1_n
rlabel polysilicon 33 0 35 36 5 S1
rlabel metal1 -58 73 -42 77 1 Vdd
rlabel metal1 -58 28 -42 32 5 GND
<< end >>
