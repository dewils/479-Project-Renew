magic
tech scmos
timestamp 1428868416
<< pwell >>
rect -1 3 27 22
<< nwell >>
rect -1 22 27 49
<< polysilicon >>
rect 4 41 6 62
rect 20 41 22 62
rect 4 24 6 33
rect 20 32 22 33
rect 20 30 30 32
rect 4 22 22 24
rect 4 15 6 17
rect 20 15 22 22
rect 4 2 6 11
rect 20 9 22 11
rect 28 2 30 30
rect 4 0 30 2
<< ndiffusion >>
rect 3 11 4 15
rect 6 11 7 15
rect 19 11 20 15
rect 22 11 23 15
<< pdiffusion >>
rect 3 33 4 41
rect 6 33 7 41
rect 19 33 20 41
rect 22 33 23 41
<< metal1 >>
rect -15 67 -12 77
rect -15 -23 -12 63
rect -8 19 -5 77
rect 38 70 41 77
rect 19 66 23 67
rect 7 62 8 66
rect -1 49 3 55
rect 23 49 27 55
rect -1 45 11 49
rect 15 45 27 49
rect -1 27 2 33
rect 8 29 11 33
rect -1 15 2 23
rect 8 15 11 25
rect 15 20 18 33
rect 24 29 27 33
rect 15 15 18 16
rect 24 15 27 25
rect -1 3 11 7
rect 15 3 27 7
rect -1 -1 3 3
rect 23 -1 27 3
rect 31 -9 34 25
rect -8 -23 -5 -13
rect 38 -23 41 66
<< metal2 >>
rect 23 67 37 70
rect -11 63 8 66
rect -19 55 -1 59
rect 27 55 45 59
rect -19 23 -1 26
rect 11 26 23 29
rect 27 26 31 29
rect 35 26 45 29
rect -5 16 14 19
rect -19 -5 -1 -1
rect 27 -5 45 -1
rect -4 -12 30 -9
<< ntransistor >>
rect 4 11 6 15
rect 20 11 22 15
<< ptransistor >>
rect 4 33 6 41
rect 20 33 22 41
<< polycontact >>
rect 3 62 7 66
rect 19 62 23 66
<< ndcontact >>
rect -1 11 3 15
rect 7 11 11 15
rect 15 11 19 15
rect 23 11 27 15
<< pdcontact >>
rect -1 33 3 41
rect 7 33 11 41
rect 15 33 19 41
rect 23 33 27 41
<< m2contact >>
rect -15 63 -11 67
rect 19 67 23 71
rect 37 66 41 70
rect 8 62 12 66
rect -1 55 3 59
rect 23 55 27 59
rect -9 15 -5 19
rect -1 23 3 27
rect 7 25 11 29
rect 23 25 27 29
rect 14 16 18 20
rect 31 25 35 29
rect -1 -5 3 -1
rect 23 -5 27 -1
rect -8 -13 -4 -9
rect 30 -13 34 -9
<< psubstratepcontact >>
rect 11 3 15 7
<< nsubstratencontact >>
rect 11 45 15 49
<< labels >>
rlabel metal2 -19 55 -1 59 7 Vdd
rlabel metal2 -19 -5 -1 -1 7 GND
rlabel metal2 -19 23 -1 26 7 A
rlabel metal2 27 55 45 59 3 Vdd
rlabel metal2 35 26 45 29 3 B
rlabel metal2 27 -5 45 -1 3 GND
rlabel metal1 -15 67 -12 77 1 shift
rlabel metal1 38 70 41 77 1 shift_n
rlabel metal1 -15 -23 -12 63 5 shift
rlabel metal1 -8 -23 -5 -13 5 B
rlabel metal1 38 -23 41 66 5 shift_n
rlabel metal1 -8 19 -5 77 1 inbit
<< end >>
