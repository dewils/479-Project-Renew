magic
tech scmos
timestamp 1428699586
<< pwell >>
rect 2 18 14 35
<< nwell >>
rect 2 35 14 56
<< polysilicon >>
rect 7 48 9 64
rect 7 30 9 40
rect 7 10 9 26
<< ndiffusion >>
rect 6 26 7 30
rect 9 26 10 30
<< pdiffusion >>
rect 6 40 7 48
rect 9 40 10 48
<< metal1 >>
rect 2 52 10 56
rect 2 48 6 52
rect 11 37 14 40
rect 11 30 14 33
rect 2 22 6 26
rect 2 18 10 22
<< metal2 >>
rect -2 56 2 60
rect 6 56 18 60
rect 15 33 18 36
rect -2 14 2 18
rect 6 14 18 18
<< ntransistor >>
rect 7 26 9 30
<< ptransistor >>
rect 7 40 9 48
<< ndcontact >>
rect 2 26 6 30
rect 10 26 14 30
<< pdcontact >>
rect 2 40 6 48
rect 10 40 14 48
<< m2contact >>
rect 2 56 6 60
rect 11 33 15 37
rect 2 14 6 18
<< psubstratepcontact >>
rect 10 18 14 22
<< nsubstratencontact >>
rect 10 52 14 56
<< labels >>
rlabel metal2 -2 56 2 60 7 Vdd
rlabel metal2 -2 14 2 18 7 GND
rlabel metal2 6 56 18 60 3 Vdd
rlabel metal2 6 14 18 18 3 GND
rlabel metal2 15 33 18 36 3 Out
rlabel polysilicon 7 48 9 64 1 In
rlabel polysilicon 7 10 9 26 5 In
<< end >>
