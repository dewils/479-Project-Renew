magic
tech scmos
timestamp 1428913770
<< pwell >>
rect 11 -9 47 8
<< nwell >>
rect 11 8 47 29
<< polysilicon >>
rect 16 21 18 33
rect 24 21 26 33
rect 40 21 42 33
rect 16 3 18 13
rect 24 3 26 13
rect 40 3 42 13
rect 48 10 50 33
rect 16 -13 18 -1
rect 24 -13 26 -1
rect 40 -13 42 -1
rect 48 -13 50 6
<< ndiffusion >>
rect 15 -1 16 3
rect 18 -1 19 3
rect 23 -1 24 3
rect 26 -1 27 3
rect 39 -1 40 3
rect 42 -1 43 3
<< pdiffusion >>
rect 15 13 16 21
rect 18 13 24 21
rect 26 13 27 21
rect 39 13 40 21
rect 42 13 43 21
<< metal1 >>
rect 7 25 19 29
rect 23 25 31 29
rect 35 25 55 29
rect 11 21 15 25
rect 35 21 39 25
rect 27 10 31 13
rect 19 6 36 10
rect 19 3 23 6
rect 43 3 47 13
rect 11 -5 15 -1
rect 27 -5 31 -1
rect 35 -5 39 -1
rect 7 -9 19 -5
rect 23 -9 31 -5
rect 35 -9 55 -5
<< ntransistor >>
rect 16 -1 18 3
rect 24 -1 26 3
rect 40 -1 42 3
<< ptransistor >>
rect 16 13 18 21
rect 24 13 26 21
rect 40 13 42 21
<< polycontact >>
rect 36 6 40 10
rect 47 6 51 10
<< ndcontact >>
rect 11 -1 15 3
rect 19 -1 23 3
rect 27 -1 31 3
rect 35 -1 39 3
rect 43 -1 47 3
<< pdcontact >>
rect 11 13 15 21
rect 27 13 31 21
rect 35 13 39 21
rect 43 13 47 21
<< psubstratepcontact >>
rect 19 -9 23 -5
rect 31 -9 35 -5
<< nsubstratencontact >>
rect 19 25 23 29
rect 31 25 35 29
<< end >>
