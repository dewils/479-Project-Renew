magic
tech scmos
timestamp 1428790139
<< pwell >>
rect 4 -14 41 8
<< nwell >>
rect 4 8 41 35
<< polysilicon >>
rect 9 27 11 48
rect 17 27 19 48
rect 33 27 35 29
rect 9 -2 11 19
rect 17 -2 19 19
rect 33 16 35 19
rect 33 -2 35 2
rect 9 -26 11 -6
rect 17 -26 19 -6
rect 33 -8 35 -6
<< ndiffusion >>
rect 8 -6 9 -2
rect 11 -6 17 -2
rect 19 -6 20 -2
rect 32 -6 33 -2
rect 35 -6 37 -2
<< pdiffusion >>
rect 8 19 9 27
rect 11 19 12 27
rect 16 19 17 27
rect 19 19 20 27
rect 32 19 33 27
rect 35 19 37 27
<< metal1 >>
rect 4 35 8 39
rect 37 35 41 39
rect 4 31 12 35
rect 16 31 28 35
rect 32 31 41 35
rect 4 27 8 31
rect 20 27 24 31
rect 28 27 32 31
rect 13 10 16 19
rect 31 11 34 12
rect 21 -2 24 6
rect 31 6 34 7
rect 38 11 41 19
rect 38 -2 41 7
rect 4 -10 8 -6
rect 28 -10 32 -6
rect 4 -14 12 -10
rect 16 -14 28 -10
rect 32 -14 41 -10
rect 4 -18 8 -14
rect 37 -18 41 -14
<< metal2 >>
rect -4 39 4 43
rect 41 39 49 43
rect 16 7 20 10
rect 24 7 30 10
rect 42 7 49 10
rect -4 -22 4 -18
rect 41 -22 49 -18
<< ntransistor >>
rect 9 -6 11 -2
rect 17 -6 19 -2
rect 33 -6 35 -2
<< ptransistor >>
rect 9 19 11 27
rect 17 19 19 27
rect 33 19 35 27
<< polycontact >>
rect 31 12 35 16
rect 31 2 35 6
<< ndcontact >>
rect 4 -6 8 -2
rect 20 -6 24 -2
rect 28 -6 32 -2
rect 37 -6 41 -2
<< pdcontact >>
rect 4 19 8 27
rect 12 19 16 27
rect 20 19 24 27
rect 28 19 32 27
rect 37 19 41 27
<< m2contact >>
rect 4 39 8 43
rect 37 39 41 43
rect 12 6 16 10
rect 20 6 24 10
rect 30 7 34 11
rect 38 7 42 11
rect 4 -22 8 -18
rect 37 -22 41 -18
<< psubstratepcontact >>
rect 12 -14 16 -10
rect 28 -14 32 -10
<< nsubstratencontact >>
rect 12 31 16 35
rect 28 31 32 35
<< end >>
