magic
tech scmos
timestamp 1428813145
<< polysilicon >>
rect 464 1600 466 1614
rect 533 1600 535 1614
rect 597 1600 599 1614
rect 663 1602 665 1614
rect 663 1600 787 1602
rect 26 800 52 802
rect 105 802 107 814
rect 56 800 150 802
rect 196 800 419 802
<< metal1 >>
rect -16 1622 -12 1694
rect -16 1522 -12 1618
rect -16 1422 -12 1518
rect -16 1322 -12 1418
rect -16 1222 -12 1318
rect -16 1122 -12 1218
rect -16 1022 -12 1118
rect -16 922 -12 1018
rect -16 822 -12 918
rect -16 722 -12 818
rect -16 622 -12 718
rect -16 522 -12 618
rect -16 422 -12 518
rect -16 322 -12 418
rect -16 222 -12 318
rect -16 122 -12 218
rect -16 52 -12 118
rect -16 22 -12 48
rect -16 -4 -12 18
rect -4 1682 0 1694
rect -4 1582 0 1678
rect -4 1482 0 1578
rect -4 1382 0 1478
rect -4 1282 0 1378
rect -4 1182 0 1278
rect -4 1082 0 1178
rect -4 982 0 1078
rect -4 882 0 978
rect 12 891 15 1694
rect 21 891 24 1694
rect -4 782 0 878
rect 53 804 56 846
rect 69 807 72 1694
rect 69 800 72 803
rect 85 800 88 845
rect 127 800 130 803
rect 192 804 195 1694
rect 463 1690 466 1694
rect 532 1690 535 1694
rect 476 1600 479 1645
rect 545 1600 548 1645
rect 585 1600 588 1694
rect 597 1690 600 1694
rect 663 1690 666 1694
rect 609 1600 612 1645
rect 706 1607 709 1694
rect 706 1600 709 1603
rect 722 1600 725 1645
rect 826 1622 830 1694
rect 764 1600 767 1603
rect 826 1522 830 1618
rect 826 1422 830 1518
rect 826 1322 830 1418
rect 826 1222 830 1318
rect 826 1122 830 1218
rect 826 1022 830 1118
rect 826 922 830 1018
rect 826 822 830 918
rect -4 682 0 778
rect -4 582 0 678
rect -4 482 0 578
rect -4 382 0 478
rect -4 282 0 378
rect -4 182 0 278
rect -4 82 0 178
rect -4 -4 0 78
rect 826 722 830 818
rect 826 622 830 718
rect 826 522 830 618
rect 826 422 830 518
rect 826 322 830 418
rect 826 222 830 318
rect 826 122 830 218
rect 826 22 830 118
rect 826 -4 830 18
rect 838 1682 842 1694
rect 838 1582 842 1678
rect 838 1482 842 1578
rect 838 1382 842 1478
rect 838 1282 842 1378
rect 838 1182 842 1278
rect 838 1082 842 1178
rect 838 982 842 1078
rect 838 882 842 978
rect 838 782 842 878
rect 838 682 842 778
rect 838 582 842 678
rect 838 482 842 578
rect 838 382 842 478
rect 838 282 842 378
rect 838 182 842 278
rect 838 82 842 178
rect 838 -4 842 78
<< metal2 >>
rect 0 1678 455 1682
rect 475 1678 524 1682
rect 544 1678 588 1682
rect 608 1678 654 1682
rect 674 1678 838 1682
rect 674 1646 721 1649
rect -12 1618 455 1622
rect 475 1618 524 1622
rect 544 1618 588 1622
rect 608 1618 654 1622
rect 674 1618 826 1622
rect 710 1604 763 1607
rect 0 1578 442 1582
rect 825 1578 838 1582
rect 825 1545 851 1548
rect -12 1518 442 1522
rect 825 1518 826 1522
rect -24 1511 442 1514
rect 0 1478 442 1482
rect 825 1478 838 1482
rect 825 1445 851 1448
rect -12 1418 442 1422
rect 825 1418 826 1422
rect -24 1411 442 1414
rect 0 1378 442 1382
rect 825 1378 838 1382
rect 825 1345 850 1348
rect -12 1318 442 1322
rect 825 1318 826 1322
rect -24 1311 442 1314
rect 0 1278 442 1282
rect 825 1278 838 1282
rect 825 1245 851 1248
rect -12 1218 442 1222
rect 825 1218 826 1222
rect -24 1211 442 1214
rect 0 1178 442 1182
rect 825 1178 838 1182
rect 825 1145 850 1148
rect -12 1118 442 1122
rect 825 1118 826 1122
rect -24 1111 442 1114
rect 0 1078 442 1082
rect 825 1078 838 1082
rect 825 1045 851 1048
rect -12 1018 442 1022
rect 825 1018 826 1022
rect -24 1011 442 1014
rect 0 978 442 982
rect 825 978 838 982
rect 825 945 850 948
rect -12 918 442 922
rect 825 918 826 922
rect -24 911 442 914
rect 53 878 96 882
rect 116 878 442 882
rect 825 878 838 882
rect 89 846 115 849
rect 825 845 851 848
rect -12 818 0 822
rect 53 818 96 822
rect 116 818 442 822
rect 825 818 826 822
rect -24 811 442 814
rect 73 804 126 807
rect 826 778 838 782
rect -24 749 0 752
rect -12 718 0 722
rect 826 678 838 682
rect -24 649 0 652
rect 826 645 851 648
rect -12 618 0 622
rect 826 578 838 582
rect -24 549 0 552
rect 826 545 851 548
rect -12 518 0 522
rect 826 478 838 482
rect -24 449 0 452
rect 826 445 851 448
rect -12 418 0 422
rect 826 378 838 382
rect -24 349 0 352
rect 826 345 851 348
rect -12 318 0 322
rect 825 278 838 282
rect -24 249 0 252
rect 826 245 851 248
rect -12 218 0 222
rect 826 178 838 182
rect -24 149 0 152
rect 826 145 851 148
rect -12 118 0 122
rect 823 78 838 82
rect -12 49 0 52
rect 826 45 851 48
rect -12 18 0 22
<< polycontact >>
rect 463 1686 467 1690
rect 532 1686 536 1690
rect 596 1686 600 1690
rect 662 1686 666 1690
rect 479 1600 483 1604
rect 548 1600 552 1604
rect 612 1600 616 1604
rect 12 887 16 891
rect 20 887 24 891
rect 52 800 56 804
rect 192 800 196 804
<< m2contact >>
rect -16 1618 -12 1622
rect -16 1518 -12 1522
rect -16 1418 -12 1422
rect -16 1318 -12 1322
rect -16 1218 -12 1222
rect -16 1118 -12 1122
rect -16 1018 -12 1022
rect -16 918 -12 922
rect -16 818 -12 822
rect -16 718 -12 722
rect -16 618 -12 622
rect -16 518 -12 522
rect -16 418 -12 422
rect -16 318 -12 322
rect -16 218 -12 222
rect -16 118 -12 122
rect -16 48 -12 52
rect -16 18 -12 22
rect -4 1678 0 1682
rect -4 1578 0 1582
rect -4 1478 0 1482
rect -4 1378 0 1382
rect -4 1278 0 1282
rect -4 1178 0 1182
rect -4 1078 0 1082
rect -4 978 0 982
rect -4 878 0 882
rect 53 846 57 850
rect 85 845 89 849
rect 69 803 73 807
rect 126 803 130 807
rect 475 1645 479 1649
rect 544 1645 548 1649
rect 608 1645 612 1649
rect 721 1645 725 1649
rect 706 1603 710 1607
rect 826 1618 830 1622
rect 763 1603 767 1607
rect 826 1518 830 1522
rect 826 1418 830 1422
rect 826 1318 830 1322
rect 826 1218 830 1222
rect 826 1118 830 1122
rect 826 1018 830 1022
rect 826 918 830 922
rect 826 818 830 822
rect -4 778 0 782
rect -4 678 0 682
rect -4 578 0 582
rect -4 478 0 482
rect -4 378 0 382
rect -4 278 0 282
rect -4 178 0 182
rect -4 78 0 82
rect 826 718 830 722
rect 826 618 830 622
rect 826 518 830 522
rect 826 418 830 422
rect 826 318 830 322
rect 826 218 830 222
rect 826 118 830 122
rect 826 18 830 22
rect 838 1678 842 1682
rect 838 1578 842 1582
rect 838 1478 842 1482
rect 838 1378 842 1382
rect 838 1278 842 1282
rect 838 1178 842 1182
rect 838 1078 842 1082
rect 838 978 842 982
rect 838 878 842 882
rect 838 778 842 782
rect 838 678 842 682
rect 838 578 842 582
rect 838 478 842 482
rect 838 378 842 382
rect 838 278 842 282
rect 838 178 842 182
rect 838 78 842 82
use ../cells/inverter1  inverter1_1
timestamp 1428803835
transform 1 0 457 0 1 1613
box -2 1 18 73
use ../cells/inverter1  inverter1_2
timestamp 1428803835
transform 1 0 526 0 1 1613
box -2 1 18 73
use ../cells/inverter1  inverter1_3
timestamp 1428803835
transform 1 0 590 0 1 1613
box -2 1 18 73
use ../cells/inverter1  inverter1_4
timestamp 1428803835
transform 1 0 656 0 1 1613
box -2 1 18 73
use ../cells/and1  and1_0
timestamp 1428803059
transform 1 0 4 0 1 839
box -4 -25 49 48
use ../cells/inverter1  inverter1_0
timestamp 1428803835
transform 1 0 98 0 1 813
box -2 1 18 73
use dbitlow  dbitlow_0
array 0 0 383 0 7 100
timestamp 1428735392
transform 1 0 442 0 1 800
box 0 0 383 100
use dbithigh  dbithigh_0
array 0 0 826 0 7 100
timestamp 1428736540
transform 1 0 0 0 1 -37
box 0 37 826 137
<< labels >>
rlabel metal1 -16 -4 -12 18 5 GND
rlabel metal1 -4 -4 0 78 5 Vdd
rlabel metal1 826 -4 830 18 5 GND
rlabel metal1 838 -4 842 78 5 Vdd
rlabel space -24 149 5 152 7 divisorin6
rlabel space -24 249 5 252 7 divisorin5
rlabel space -24 349 5 352 7 divisorin4
rlabel space -24 449 5 452 7 divisorin3
rlabel space -24 549 5 552 7 divisorin2
rlabel space -24 649 5 652 7 divisorin1
rlabel space -24 749 5 752 7 divisorin0
rlabel space -24 811 445 814 7 dividenin7
rlabel space -24 911 445 914 7 dividenin6
rlabel space -24 1011 445 1014 7 dividenin5
rlabel space -24 1111 445 1114 7 dividenin4
rlabel space -24 1211 445 1214 7 dividenin3
rlabel space -24 1311 445 1314 7 dividenin2
rlabel space -24 1411 445 1414 7 dividenin1
rlabel space -24 1511 445 1514 7 dividenin0
rlabel metal1 -16 1622 -12 1694 1 GND
rlabel metal1 -4 1682 0 1694 1 Vdd
rlabel metal1 12 891 15 1694 1 clk
rlabel metal1 21 891 24 1694 1 load
rlabel metal1 69 807 72 1694 1 reset_n
rlabel metal1 192 804 195 1694 1 add_n
rlabel metal1 463 1690 466 1694 1 sel0
rlabel metal1 532 1690 535 1694 1 sel1
rlabel space 585 1555 588 1694 1 inbit
rlabel metal1 597 1690 600 1694 1 shift
rlabel metal1 663 1690 666 1694 1 clk
rlabel metal1 706 1607 709 1694 1 reset_n
rlabel metal1 838 1682 842 1694 1 Vdd
rlabel metal1 826 1622 830 1694 1 GND
rlabel space 822 45 851 48 3 remainder6
rlabel space 822 145 851 148 3 remainder5
rlabel space 822 245 851 248 3 remainder4
rlabel space 822 345 851 348 3 remainder3
rlabel space 822 445 851 448 3 remainder2
rlabel space 822 545 851 548 3 remainder1
rlabel space 822 645 851 648 3 remainder0
rlabel space 822 845 851 848 3 quotient7
rlabel space 822 945 850 948 3 quotient6
rlabel space 822 1045 851 1048 3 quotient5
rlabel space 822 1145 850 1148 3 quotient4
rlabel space 822 1245 851 1248 3 quotient3
rlabel space 822 1345 850 1348 3 quotient2
rlabel space 822 1445 851 1448 3 quotient1
rlabel space 822 1545 851 1548 3 quotient0
<< end >>
