magic
tech scmos
timestamp 1428701418
<< pwell >>
rect -1 3 27 22
<< nwell >>
rect -1 22 27 49
<< polysilicon >>
rect 4 41 6 77
rect 20 44 22 77
rect 20 42 31 44
rect 20 41 22 42
rect 4 27 6 33
rect 20 31 22 33
rect 4 25 22 27
rect 4 15 6 17
rect 20 15 22 25
rect 4 -5 6 11
rect 20 -14 22 11
rect 4 -16 22 -14
rect 4 -23 6 -16
rect 20 -20 25 -18
rect 29 -20 31 42
rect 20 -23 22 -20
<< ndiffusion >>
rect 3 11 4 15
rect 6 11 7 15
rect 19 11 20 15
rect 22 11 23 15
<< pdiffusion >>
rect 3 33 4 41
rect 6 33 7 41
rect 19 33 20 41
rect 22 33 23 41
<< metal1 >>
rect -8 32 -5 77
rect -1 49 3 55
rect 23 49 27 55
rect -1 45 11 49
rect 15 45 27 49
rect -1 22 2 33
rect -1 15 2 18
rect 8 22 11 33
rect 15 32 18 33
rect 8 15 11 18
rect 15 15 18 28
rect 24 22 27 33
rect 24 15 27 18
rect 33 7 36 18
rect -1 3 11 7
rect 15 3 27 7
rect -8 -23 -5 3
rect -1 -1 3 3
rect 23 -1 27 3
rect 7 -9 10 -5
rect 25 -16 28 -13
<< metal2 >>
rect -12 55 -1 59
rect 27 55 40 59
rect -4 28 14 31
rect -12 18 -2 21
rect 12 18 24 21
rect 28 18 32 21
rect 36 18 40 21
rect -4 3 33 6
rect -12 -5 -1 -1
rect 27 -5 40 -1
rect 11 -13 24 -10
<< ntransistor >>
rect 4 11 6 15
rect 20 11 22 15
<< ptransistor >>
rect 4 33 6 41
rect 20 33 22 41
<< polycontact >>
rect 6 -5 10 -1
rect 25 -20 29 -16
<< ndcontact >>
rect -1 11 3 15
rect 7 11 11 15
rect 15 11 19 15
rect 23 11 27 15
<< pdcontact >>
rect -1 33 3 41
rect 7 33 11 41
rect 15 33 19 41
rect 23 33 27 41
<< m2contact >>
rect -1 55 3 59
rect 23 55 27 59
rect -8 28 -4 32
rect -2 18 2 22
rect 14 28 18 32
rect 8 18 12 22
rect 24 18 28 22
rect 32 18 36 22
rect -8 3 -4 7
rect 33 3 37 7
rect -1 -5 3 -1
rect 23 -5 27 -1
rect 7 -13 11 -9
rect 24 -13 28 -9
<< psubstratepcontact >>
rect 11 3 15 7
<< nsubstratencontact >>
rect 11 45 15 49
<< labels >>
rlabel polysilicon 4 41 6 77 1 shift
rlabel polysilicon 20 41 22 77 1 noshift
rlabel metal2 -12 55 -1 59 7 Vdd
rlabel metal2 27 55 40 59 3 Vdd
rlabel metal2 -12 -5 -1 -1 7 GND
rlabel metal2 27 -5 40 -1 3 GND
rlabel polysilicon 4 -23 6 -14 5 shift
rlabel polysilicon 20 -23 22 -18 5 noshift
rlabel metal1 -8 -23 -5 3 5 B
rlabel metal2 36 18 40 21 3 B
rlabel metal2 -12 18 -2 21 7 A
rlabel metal1 -8 32 -5 77 1 inbit
<< end >>
