magic
tech scmos
timestamp 1428736404
<< pwell >>
rect -109 26 137 58
<< nwell >>
rect -109 58 137 90
<< polysilicon >>
rect -104 82 -102 108
rect 120 102 122 108
rect -17 100 122 102
rect -82 82 -80 84
rect -60 82 -58 84
rect -41 82 -39 84
rect -33 82 -31 93
rect -17 82 -15 100
rect -1 82 1 84
rect 4 82 6 93
rect 20 82 22 84
rect 37 82 39 84
rect 45 82 47 93
rect 61 82 63 100
rect 81 82 83 84
rect 98 82 100 84
rect 104 82 106 93
rect 110 82 112 100
rect 129 82 131 84
rect -104 60 -102 72
rect -82 71 -80 72
rect -104 58 -91 60
rect -60 60 -58 72
rect -87 58 -58 60
rect -104 39 -102 58
rect -82 39 -80 40
rect -60 39 -58 40
rect -41 39 -39 72
rect -33 61 -31 72
rect -33 59 -28 61
rect -33 39 -31 59
rect -17 39 -15 72
rect -1 39 1 72
rect 4 39 6 72
rect 20 69 22 72
rect 20 39 22 42
rect 37 39 39 72
rect 45 39 47 72
rect 61 39 63 72
rect 81 69 83 72
rect 81 39 83 42
rect 98 39 100 72
rect 104 39 106 72
rect 110 39 112 72
rect 129 69 131 72
rect -104 8 -102 34
rect -82 32 -80 34
rect -60 32 -58 34
rect -41 25 -39 34
rect -33 32 -31 34
rect -17 32 -15 34
rect -1 25 1 34
rect 4 32 6 34
rect 20 32 22 34
rect 37 25 39 34
rect 45 32 47 34
rect 61 32 63 34
rect 81 32 83 34
rect 98 25 100 34
rect 104 32 106 34
rect 110 32 112 34
rect -41 23 100 25
rect 120 8 122 42
rect 129 39 131 42
rect 129 32 131 34
<< ndiffusion >>
rect -105 34 -104 39
rect -102 34 -98 39
rect -86 34 -82 39
rect -80 34 -76 39
rect -64 34 -60 39
rect -58 34 -54 39
rect -42 34 -41 39
rect -39 34 -38 39
rect -34 34 -33 39
rect -31 34 -30 39
rect -18 34 -17 39
rect -15 34 -14 39
rect -2 34 -1 39
rect 1 34 4 39
rect 6 34 7 39
rect 19 34 20 39
rect 22 34 24 39
rect 36 34 37 39
rect 39 34 40 39
rect 44 34 45 39
rect 47 34 48 39
rect 60 34 61 39
rect 63 34 64 39
rect 76 34 81 39
rect 83 34 85 39
rect 97 34 98 39
rect 100 34 104 39
rect 106 34 110 39
rect 112 34 113 39
rect 128 34 129 39
rect 131 34 133 39
<< pdiffusion >>
rect -105 72 -104 82
rect -102 72 -98 82
rect -86 72 -82 82
rect -80 72 -76 82
rect -64 72 -60 82
rect -58 72 -54 82
rect -42 72 -41 82
rect -39 72 -38 82
rect -34 72 -33 82
rect -31 72 -30 82
rect -18 72 -17 82
rect -15 72 -14 82
rect -2 72 -1 82
rect 1 72 4 82
rect 6 72 7 82
rect 19 72 20 82
rect 22 72 24 82
rect 36 72 37 82
rect 39 72 40 82
rect 44 72 45 82
rect 47 72 48 82
rect 60 72 61 82
rect 63 72 64 82
rect 76 72 81 82
rect 83 72 85 82
rect 97 72 98 82
rect 100 72 104 82
rect 106 72 110 82
rect 112 72 113 82
rect 128 72 129 82
rect 131 72 133 82
<< metal1 >>
rect -33 97 -30 103
rect 4 97 7 103
rect 45 97 48 103
rect 103 97 106 103
rect -105 86 -94 90
rect -90 86 -72 90
rect -68 86 -54 90
rect -50 86 -38 90
rect -34 86 -26 90
rect -22 86 -10 90
rect -6 86 11 90
rect 15 86 28 90
rect 32 86 40 90
rect 44 86 52 90
rect 56 86 72 90
rect 76 86 85 90
rect 89 86 120 90
rect 124 86 133 90
rect -109 82 -105 86
rect -46 82 -42 86
rect -30 82 -26 86
rect -6 82 -2 86
rect 15 82 19 86
rect 32 82 36 86
rect 48 82 52 86
rect 64 82 68 86
rect 93 82 97 86
rect 124 82 128 86
rect -97 48 -94 72
rect -90 62 -87 72
rect -83 65 -80 67
rect -83 56 -80 61
rect -75 57 -72 72
rect -97 39 -94 44
rect -83 44 -80 52
rect -90 39 -87 44
rect -75 39 -72 53
rect -68 56 -65 72
rect -53 65 -50 72
rect -38 69 -35 72
rect -22 69 -19 72
rect -68 39 -65 52
rect -60 44 -57 45
rect -53 39 -50 61
rect -28 55 -25 58
rect -13 54 -10 72
rect 8 61 11 72
rect 8 53 11 57
rect 18 54 21 65
rect -38 39 -35 42
rect -22 39 -19 42
rect -13 39 -10 50
rect 8 39 11 49
rect 18 46 21 50
rect 25 54 28 72
rect 40 69 43 72
rect 56 69 59 72
rect 72 69 75 72
rect 79 61 82 65
rect 25 39 28 50
rect 79 46 82 57
rect 86 64 89 72
rect 114 64 117 72
rect 127 64 130 65
rect 40 39 43 42
rect 56 39 59 42
rect 72 39 75 42
rect 86 39 89 60
rect 114 39 117 60
rect 120 46 123 50
rect 127 46 130 60
rect 134 60 137 72
rect 134 39 137 56
rect -109 30 -105 34
rect -46 30 -42 34
rect -30 30 -26 34
rect -6 30 -2 34
rect 15 30 19 34
rect 32 30 36 34
rect 48 30 52 34
rect 64 30 68 34
rect 93 30 97 34
rect 124 30 128 34
rect -105 26 -94 30
rect -90 26 -72 30
rect -68 26 -54 30
rect -50 26 -38 30
rect -34 26 -26 30
rect -22 26 -11 30
rect -7 26 11 30
rect 15 26 27 30
rect 31 26 40 30
rect 44 26 52 30
rect 56 26 72 30
rect 76 26 85 30
rect 89 26 113 30
rect 117 26 133 30
rect -41 16 -38 19
<< metal2 >>
rect -29 104 4 107
rect 8 104 45 107
rect 49 104 103 107
rect -113 86 -109 90
rect 137 86 141 90
rect -34 65 -23 68
rect 44 65 56 68
rect 60 65 72 68
rect -80 62 -54 65
rect 11 58 78 61
rect 90 60 113 63
rect 117 60 126 63
rect -113 53 -84 56
rect 138 57 141 60
rect -72 53 -68 56
rect -64 55 -24 56
rect -64 53 -28 55
rect -10 50 7 53
rect 11 50 17 53
rect 29 50 120 53
rect -94 45 -90 48
rect -86 45 -60 48
rect -34 43 -23 46
rect 44 42 56 45
rect 60 42 72 45
rect -113 26 -109 30
rect 137 26 141 30
rect -113 12 -42 15
rect -38 12 141 15
<< ntransistor >>
rect -104 34 -102 39
rect -82 34 -80 39
rect -60 34 -58 39
rect -41 34 -39 39
rect -33 34 -31 39
rect -17 34 -15 39
rect -1 34 1 39
rect 4 34 6 39
rect 20 34 22 39
rect 37 34 39 39
rect 45 34 47 39
rect 61 34 63 39
rect 81 34 83 39
rect 98 34 100 39
rect 104 34 106 39
rect 110 34 112 39
rect 129 34 131 39
<< ptransistor >>
rect -104 72 -102 82
rect -82 72 -80 82
rect -60 72 -58 82
rect -41 72 -39 82
rect -33 72 -31 82
rect -17 72 -15 82
rect -1 72 1 82
rect 4 72 6 82
rect 20 72 22 82
rect 37 72 39 82
rect 45 72 47 82
rect 61 72 63 82
rect 81 72 83 82
rect 98 72 100 82
rect 104 72 106 82
rect 110 72 112 82
rect 129 72 131 82
<< polycontact >>
rect -33 93 -29 97
rect 4 93 8 97
rect 45 93 49 97
rect 103 93 107 97
rect -83 67 -79 71
rect -91 58 -87 62
rect -83 40 -79 44
rect -61 40 -57 44
rect -28 58 -24 62
rect 18 65 22 69
rect 18 42 22 46
rect 79 65 83 69
rect 79 42 83 46
rect 127 65 131 69
rect 120 42 124 46
rect 127 42 131 46
rect -42 19 -38 23
<< ndcontact >>
rect -109 34 -105 39
rect -98 34 -94 39
rect -90 34 -86 39
rect -76 34 -72 39
rect -68 34 -64 39
rect -54 34 -50 39
rect -46 34 -42 39
rect -38 34 -34 39
rect -30 34 -26 39
rect -22 34 -18 39
rect -14 34 -10 39
rect -6 34 -2 39
rect 7 34 11 39
rect 15 34 19 39
rect 24 34 28 39
rect 32 34 36 39
rect 40 34 44 39
rect 48 34 52 39
rect 56 34 60 39
rect 64 34 68 39
rect 72 34 76 39
rect 85 34 89 39
rect 93 34 97 39
rect 113 34 117 39
rect 124 34 128 39
rect 133 34 137 39
<< pdcontact >>
rect -109 72 -105 82
rect -98 72 -94 82
rect -90 72 -86 82
rect -76 72 -72 82
rect -68 72 -64 82
rect -54 72 -50 82
rect -46 72 -42 82
rect -38 72 -34 82
rect -30 72 -26 82
rect -22 72 -18 82
rect -14 72 -10 82
rect -6 72 -2 82
rect 7 72 11 82
rect 15 72 19 82
rect 24 72 28 82
rect 32 72 36 82
rect 40 72 44 82
rect 48 72 52 82
rect 56 72 60 82
rect 64 72 68 82
rect 72 72 76 82
rect 85 72 89 82
rect 93 72 97 82
rect 113 72 117 82
rect 124 72 128 82
rect 133 72 137 82
<< m2contact >>
rect -33 103 -29 107
rect 4 103 8 107
rect 45 103 49 107
rect 103 103 107 107
rect -109 86 -105 90
rect 133 86 137 90
rect -84 61 -80 65
rect -84 52 -80 56
rect -76 53 -72 57
rect -98 44 -94 48
rect -90 44 -86 48
rect -38 65 -34 69
rect -23 65 -19 69
rect -54 61 -50 65
rect -68 52 -64 56
rect -60 45 -56 49
rect -28 51 -24 55
rect 7 57 11 61
rect -14 50 -10 54
rect -38 42 -34 46
rect -23 42 -19 46
rect 7 49 11 53
rect 17 50 21 54
rect 40 65 44 69
rect 56 65 60 69
rect 72 65 76 69
rect 78 57 82 61
rect 25 50 29 54
rect 86 60 90 64
rect 113 60 117 64
rect 126 60 130 64
rect 40 42 44 46
rect 56 42 60 46
rect 72 42 76 46
rect 120 50 124 54
rect 134 56 138 60
rect -109 26 -105 30
rect 133 26 137 30
rect -42 12 -38 16
<< psubstratepcontact >>
rect -94 26 -90 30
rect -72 26 -68 30
rect -54 26 -50 30
rect -38 26 -34 30
rect -26 26 -22 30
rect -11 26 -7 30
rect 11 26 15 30
rect 27 26 31 30
rect 40 26 44 30
rect 52 26 56 30
rect 72 26 76 30
rect 85 26 89 30
rect 113 26 117 30
<< nsubstratencontact >>
rect -94 86 -90 90
rect -72 86 -68 90
rect -54 86 -50 90
rect -38 86 -34 90
rect -26 86 -22 90
rect -10 86 -6 90
rect 11 86 15 90
rect 28 86 32 90
rect 40 86 44 90
rect 52 86 56 90
rect 72 86 76 90
rect 85 86 89 90
rect 120 86 124 90
<< labels >>
rlabel polysilicon -104 82 -102 108 1 add_n
rlabel polysilicon -104 8 -102 34 5 add_n
rlabel metal2 -113 53 -84 56 7 B
rlabel polysilicon 120 8 122 26 5 X
rlabel polysilicon 120 100 122 108 1 C
rlabel metal2 138 57 141 60 3 Z
rlabel metal2 -113 86 -109 90 7 Vdd
rlabel metal2 -113 26 -109 30 7 GND
rlabel metal2 137 86 141 90 3 Vdd
rlabel metal2 137 26 141 30 3 GND
rlabel metal2 -113 12 -42 15 7 A
rlabel metal2 -38 12 141 15 3 A
<< end >>
