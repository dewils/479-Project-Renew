magic
tech scmos
timestamp 1428294818
<< pwell >>
rect -5 6 31 26
<< nwell >>
rect -5 26 31 49
<< polysilicon >>
rect 4 41 6 77
rect 20 41 22 77
rect 4 31 6 33
rect 20 31 22 33
rect 4 19 6 21
rect 20 19 22 21
rect 4 -23 6 15
rect 20 -23 22 15
<< ndiffusion >>
rect 3 15 4 19
rect 6 15 7 19
rect 19 15 20 19
rect 22 15 23 19
<< pdiffusion >>
rect 3 33 4 41
rect 6 33 7 41
rect 19 33 20 41
rect 22 33 23 41
<< metal1 >>
rect -5 45 11 49
rect 15 45 31 49
rect -1 32 2 33
rect -1 19 2 28
rect 8 32 11 33
rect 8 19 11 28
rect 15 24 18 33
rect 15 19 18 20
rect 24 32 27 33
rect 24 19 27 28
rect -5 6 11 10
rect 15 6 31 10
<< metal2 >>
rect -5 29 -2 32
rect 12 29 24 32
rect 28 29 31 32
rect -5 20 14 23
<< ntransistor >>
rect 4 15 6 19
rect 20 15 22 19
<< ptransistor >>
rect 4 33 6 41
rect 20 33 22 41
<< ndcontact >>
rect -1 15 3 19
rect 7 15 11 19
rect 15 15 19 19
rect 23 15 27 19
<< pdcontact >>
rect -1 33 3 41
rect 7 33 11 41
rect 15 33 19 41
rect 23 33 27 41
<< m2contact >>
rect -2 28 2 32
rect 8 28 12 32
rect 14 20 18 24
rect 24 28 28 32
<< psubstratepcontact >>
rect 11 6 15 10
<< nsubstratencontact >>
rect 11 45 15 49
<< labels >>
rlabel metal1 -5 45 11 49 1 Vdd
rlabel metal1 -5 6 11 10 5 GND
rlabel metal2 -5 29 -2 32 7 A
rlabel metal2 -5 20 14 23 7 inbit
rlabel metal2 28 29 31 32 3 B
rlabel polysilicon 4 41 6 77 1 shift
rlabel polysilicon 20 41 22 77 1 noshift
rlabel polysilicon 4 -23 6 15 5 noshift
rlabel polysilicon 20 -23 22 15 5 shift
<< end >>
